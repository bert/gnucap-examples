* Spice netlister for gnetlist
V1 2 1 DC 10V
V2 4 3 DC 5V
V3 0 3 DC 3V
R1 1 2 220
R2 2 3 4k7
R3 4 5 3k3
R4 3 5 10k
R5 0 1 22k
R6 0 5 15k
.END
