* Coilcraft XGL4020-102 1.0uH

.param L1_R1 = 34
.param L1_R2 = 8.2e-3
.param L1_C= 6.87pF
.param L1_K1 = 1e-6
.param L1_K2 = 0.236
.param L1_K3=1
.param L1_K4 = 9e-3
.param L1_K5 = 4e-3

V1 Vin 0 AC 1
R2 N001 Vin {L1_R2}
R1 0 N002 {L1_R1}
C1 N002 N001 {L1_C}
G§Rvar1 N001 0 N001 0 LAPLACE=+1/{L1_K2}/(-S*S/4/PI^2)^0.25
G§Rvar2 N001 N003 N001 N003 LAPLACE=+1/{L1_K1}/(-S*S/4/PI^2)^0.25
G§Lvar1 N003 0 N003 0 LAPLACE=+1/(S*1e-6*({L1_K3}-({L1_K4}*LOG({L1_K5}*(abs(S)/(2*pi))))))
R3 N003 0 100Meg

.ac dec 250 1e5 5e8
* NOTE: \nInd   = IM(V(Vin)/I(R2))/(2*PI*Frequency)\nImp  = V(Vin)/I(R2)\nESR= RE(V(Vin)/I(R2))
.backanno
.end
