.title eg3.ckt

I1 1 4 DC 2mA
V1 1 0 DC 5V

* begin vcvs expansion, e<name>
E1 5 2 1 3 0.4
Isense_E1 1 3 dc 0
IOut_E1 5 2 dc 0
* end vcvs expansion

* begin cccs expansion, f<name>
F1 5 6 Vsense_F1 1
Vsense_F1 R1 3e-2 dc 0
* end cccs expansion

* begin vccs expansion, g<name>
G1 2 3 4 6 1.3
IMeasure_G1 4 6 dc 0
* end vccs expansion

* begin ccvs expansion, h<name>
H1 3 0 Vsense_H1 1
Vsense_H1 R3 1 dc 0
IOut_H1 3 0 dc 0
* end ccvs expansion

R1 4 5 2.2  
R2 1 2 470  
R3 0 2 330  
R4 3 6 1k  
R5 5 6 1e4

.print dc v(2) z(2)

.dc

.end
