.TITLE PELTZ OSCILLATOR - TRANSIENT RESPONSE

.MODEL 2N3904 NPN

VEE 5 0 -5

C1 0 2 100p
L1 0 2 100u
R1 4 5 10k
R2 0 1 4.7k
R3 2 3 4.7k
Q1 2 1 4 2N3904
Q2 0 3 4 2N3904

.PRINT OP Iter(0) V(2)

.PRINT TRAN V(2) V(4)

*     FROM  TO       STEP  OPTIONS
.TRAN 0     0.00002  1e-8

.END
