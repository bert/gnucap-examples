eg4.ckt
* VOLTAGE SOURCES IN PARALLEL

V1 1 0 10.0
V2 1 0 10.2
.print dc v(1) i(V1) i(V2)
.dc
.end
